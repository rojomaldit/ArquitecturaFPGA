module imem (input logic [5:0] addr,
				 output logic [31:0] q);
			
	logic [31:0] rom [0:18] = '{
                              32'h91003c0a,
                              32'hd503201f,
                              32'hd503201f,
                              32'hd503201f,
                              32'hf800000a,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000,
                              32'h00000000
                             };


	assign q = rom[addr];
endmodule
