module signext_tb();
	logic[31:0] a;
	logic[63:0] y;
	
	signext test(a, y);
	
	initial begin
		//LDUR
		a = 32'b11111000010_000000001_00_00000_00000; #5;
		a = 32'b11111000010_100000001_00_00000_00000; #5;
		
		//STUR
		a = 32'b11111000000_000001001_00_00000_00000; #5;
		a = 32'b11111000000_100100001_00_00000_00000; #5;
		
		//CBZ
		a = 32'b10110100000_000000001_00_00000_00000; #5;
		a = 32'b10110100000_100000001_00_00000_00000; #5;
		
		//NO EXPRESION
		a = 32'b11111111111_000000001_00_00000_00000; #5;
		a = 32'b11111011001_100000001_00_00000_00000; #5;
		
	end

endmodule 